module rom (
    input [5:0]addr,
    input clk,
    output reg [7:0]q
);

always @(posedge clk) begin
    case (addr)
//    3'b000: q = 8'b01011011; // [
//    3'b001: q = 8'b01000110; // F
//    3'b010: q = 8'b01010000; // P
//    3'b011: q = 8'b01000111; // G
//    3'b100: q = 8'b01000001; // A
//    3'b101: q = 8'b01011101; // ]
//    3'b110: q = 8'b00001101; // \r
//    3'b111: q = 8'b00001010; // \n
        6'b000000: q = 8'b00100000; // ' '
        6'b000001: q = 8'b01111100; // '|'
        6'b000010: q = 8'b01011100; // '\'
        6'b000011: q = 8'b01011111; // '_'
        6'b000100: q = 8'b01011111; // '_'
        6'b000101: q = 8'b00101111; // '/'
        6'b000110: q = 8'b00101100; // ','
        6'b000111: q = 8'b01111100; // '|'
        6'b001000: q = 8'b00100000; // ' '
        6'b001001: q = 8'b00100000; // ' '
        6'b001010: q = 8'b00100000; // ' '
        6'b001011: q = 8'b00101000; // '('
        6'b001100: q = 8'b01100000; // '`'
        6'b001101: q = 8'b01011100; // '\'
        6'b001110: q = 8'b00001101; // '\r'
        6'b001111: q = 8'b00001010; // '\n'
        6'b010000: q = 8'b00100000; // ' '
        6'b010001: q = 8'b01111100; // '|'
        6'b010010: q = 8'b01011111; // '_'
        6'b010011: q = 8'b00100000; // ' '
        6'b010100: q = 8'b01011111; // '_'
        6'b010101: q = 8'b00100000; // ' '
        6'b010110: q = 8'b00100000; // ' '
        6'b010111: q = 8'b01111100; // '|'
        6'b011000: q = 8'b00101110; // '.'
        6'b011001: q = 8'b00101101; // '-'
        6'b011010: q = 8'b00101101; // '-'
        6'b011011: q = 8'b00101110; // '.'
        6'b011100: q = 8'b00101001; // ')'
        6'b011101: q = 8'b00100000; // ' '
        6'b011110: q = 8'b00101001; // ')'
        6'b011111: q = 8'b00001101; // '\r'
        6'b100000: q = 8'b00001010; // '\n'
        6'b100001: q = 8'b00100000; // ' '
        6'b100010: q = 8'b00101000; // '('
        6'b100011: q = 8'b00100000; // ' '
        6'b100100: q = 8'b01010100; // 'T'
        6'b100101: q = 8'b00100000; // ' '
        6'b100110: q = 8'b00100000; // ' '
        6'b100111: q = 8'b00100000; // ' '
        6'b101000: q = 8'b00101001; // ')'
        6'b101001: q = 8'b00100000; // ' '
        6'b101010: q = 8'b00100000; // ' '
        6'b101011: q = 8'b00100000; // ' '
        6'b101100: q = 8'b00100000; // ' '
        6'b101101: q = 8'b00100000; // ' '
        6'b101110: q = 8'b00101111; // '/'
        6'b101111: q = 8'b00001101; // '\r'
        6'b110000: q = 8'b00001010; // '\n'
        6'b110001: q = 8'b00101000; // '('
        6'b110010: q = 8'b00101000; // '('
        6'b110011: q = 8'b00101000; // '('
        6'b110100: q = 8'b01011110; // '^'
        6'b110101: q = 8'b01011111; // '_'
        6'b110110: q = 8'b00101000; // '('
        6'b110111: q = 8'b00101000; // '('
        6'b111000: q = 8'b00101000; // '('
        6'b111001: q = 8'b00101111; // '/'
        6'b111010: q = 8'b00101000; // '('
        6'b111011: q = 8'b00101000; // '('
        6'b111100: q = 8'b01011111; // '_'
        6'b111101: q = 8'b00101111; // '/'
        6'b111110: q = 8'b00001101; // '\r'
        6'b111111: q = 8'b00001010; // '\n'
    endcase
end

endmodule
